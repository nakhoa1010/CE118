library verilog;
use verilog.vl_types.all;
entity Bai1_vlg_vec_tst is
end Bai1_vlg_vec_tst;
