library verilog;
use verilog.vl_types.all;
entity Bai1_vlg_check_tst is
    port(
        O               : in     vl_logic;
        Q0              : in     vl_logic;
        Q1              : in     vl_logic;
        Q2              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Bai1_vlg_check_tst;
